--Reyes Mendoza Miriam Guadalupe
--Guerrero Prado Issac Alexander
--No. Cuenta 315569131
--No. Cuenta 317231117


library ieee;
use ieee.std_logic_1164.all;

entity divf is
port(
clk, reset, stop: in std_logic;
cuenta: out std_logic_vector(3 downto 0));
end;

architecture arq of divf is
signal clkl: std_logic;
begin
end;