library ieee;
use ieee.std_logic_1164.all;

entity divf3 is
generic(num: integer:=25000000);
port(clk: in std_logic;
	  sal: buffer std_logic);
end entity;

architecture arqdivf of divf3 is

signal conteo: integer range 0 to num;

begin
   process (clk)
   begin
      if rising_edge (clk) then
			if(conteo=num) then
				conteo<=0;
				sal<= not sal;
			else
				conteo<=conteo+1;
			end if;
      end if;
      end process;
end architecture;